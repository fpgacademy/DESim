// choose VGA resolution: Options are:
//
// `define VGA_640_480
`define VGA_320_240
//`define VGA_160_120

